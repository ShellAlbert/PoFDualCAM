`timescale 1ns/1ns


module tb_top();
// ADC Core Simulation model is not available
	
endmodule
